package adsb_decoder_p is

    constant INPUT_POWER_WIDTH  :   natural     := 32 ;

end package ;

